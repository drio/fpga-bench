`default_nettype none `timescale 1 ns / 1ns

module sha256(
  input logic clk
);

endmodule
